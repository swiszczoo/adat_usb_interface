module nrzi_phase_lock_decoder (
    input logic     clk_i,
    input logic     clk_x4_i,
    input logic     nrzi_i,
    output logic    data_o,
    output logic    valid_o
);
    // TODO: write logic
endmodule
