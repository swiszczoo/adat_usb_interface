module nrzi_encoder (
    input           data_i,
    input           clk_x4_i,
    output          data_o
);
    
endmodule
