module main;

endmodule
